`default_nettype none `timescale 1ns / 1ps

/* This testbench just instantiates the module and makes some convenient wires
   that can be driven / tested by the cocotb test.py.
*/
module tb ();

  // Dump the signals to a VCD file. You can view it with gtkwave.
  initial begin
    $dumpfile("tb.vcd");
    $dumpvars(0, tb);
    #1;
  end

  // Wire up the inputs and outputs:
  reg clk;
  reg rst_n;
  reg ena;
  reg [7:0] ui_in;
  reg [7:0] uio_in;
  wire [7:0] uo_out;
  wire [7:0] uio_out;
  wire [7:0] uio_oe;
  
  //wire for testing with cocotb
  wire reset = rst_n;
  wire [10:0] m_axis_fir_tdata; //FIR OUTPUT DATA
  wire s_set_coeffs;
  wire s_axis_fir_tvalid;
  wire [7:0] s_axis_fir_tdata; //FIR INPUT DATA 
  
  //assign inputs
  assign s_axis_fir_tdata = ui_in[7:0]; //8 Bit in
  assign s_axis_fir_tvalid = uio_in[7];
  assign s_set_coeffs = uio_in[6];
  
  //assign outputs
  assign uo_out = m_axis_fir_tdata[7:0]; //8Bits output
  assign uio_out[2:0] = m_axis_fir_tdata[10:8]; //2Bits output
  
  
  
      
  //remainder - set to defined state and config
  assign uio_oe[7:0] = 8'b00111111;
  assign uio_out[5:3] = 3'b000;
  assign uio_out[7:6] = 2'b00;

    
    

  // Replace tt_um_example with your module name:
  tt_um_haeuslermarkus_fir_filter tt_um_haeuslermarkus_fir_filter_inst (

      // Include power ports for the Gate Level test:
`ifdef GL_TEST
      .VPWR(1'b1),
      .VGND(1'b0),
`endif

      .ui_in  (ui_in),    // Dedicated inputs
      .uo_out (uo_out),   // Dedicated outputs
      .uio_in (uio_in),   // IOs: Input path
      .uio_out(uio_out),  // IOs: Output path
      .uio_oe (uio_oe),   // IOs: Enable path (active high: 0=input, 1=output)
      .ena    (ena),      // enable - goes high when design is selected
      .clk    (clk),      // clock
      .rst_n  (rst_n)     // not reset
  );

endmodule
